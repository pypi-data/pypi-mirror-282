// DESCRIPTION: Verilator: Verilog Test module
//
// This file ONLY is placed under the Creative Commons Public Domain, for
// any use, without warranty, 2023 by Antmicro Ltd.
// SPDX-License-Identifier: CC0-1.0

module t (/*AUTOARG*/);

   class Bar #(type T=int) extends T;
   endclass

   initial begin
      Bar#() bar;
      $stop;
   end
endmodule
