// DESCRIPTION: Verilator: Dotted reference that uses another dotted reference
// as the select expression
//
// This file ONLY is placed into the Public Domain, for any use,
// without warranty, 2023 by Wilson Snyder.
// SPDX-License-Identifier: CC0-1.0

`include "t/t_debug_inputs_a.v"

module t_debug_inputs (/*AUTOARG*/);
endmodule
