// DESCRIPTION: Verilog::Preproc: Example source code
// This file ONLY is placed under the Creative Commons Public Domain, for
// any use, without warranty, 2000-2011 by Wilson Snyder.
// SPDX-License-Identifier: CC0-1.0

`define T_PREPROC_INC4
