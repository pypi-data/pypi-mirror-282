// DESCRIPTION: Verilator: Verilog Test module
//
// This file ONLY is placed under the Creative Commons Public Domain, for
// any use, without warranty, 2019 by Wilson Snyder.
// SPDX-License-Identifier: CC0-1.0

// Legal with ANSI Verilog 2001 style ports
module t
  (
   output wire ok_ow,
   output reg  ok_or);

   wire ok_o_w;
   reg   ok_o_r;
endmodule
