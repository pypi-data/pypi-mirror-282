// DESCRIPTION: Verilator: Verilog Test module
//
// This file ONLY is placed under the Creative Commons Public Domain, for
// any use, without warranty, 2023 by Wilson Snyder.
// SPDX-License-Identifier: CC0-1.0

module sub;
   // verilator lint_off WIDTHTRUNC
   int warn_sub = 64'h1;  // Suppressed
endmodule
